module SM4_SBOX(
	input      [7:0]    sm4_box_in,
	output reg [7:0]    sm4_box_out													
);

always @(*) begin
	case(sm4_box_in)
		8'h00:	  sm4_box_out	<=	8'hd6;
		8'h01:	  sm4_box_out	<=	8'h90;
		8'h02:	  sm4_box_out	<=	8'he9;
		8'h03:	  sm4_box_out	<=	8'hfe;
		8'h04:	  sm4_box_out	<=	8'hcc;
		8'h05:	  sm4_box_out	<=	8'he1;
		8'h06:	  sm4_box_out	<=	8'h3d;
		8'h07:	  sm4_box_out	<=	8'hb7;
		8'h08:	  sm4_box_out	<=	8'h16;
		8'h09:	  sm4_box_out	<=	8'hb6;
		8'h0a:	  sm4_box_out	<=	8'h14;
		8'h0b:	  sm4_box_out	<=	8'hc2;
		8'h0c:	  sm4_box_out	<=	8'h28;
		8'h0d:	  sm4_box_out	<=	8'hfb;
		8'h0e:	  sm4_box_out	<=	8'h2c;
		8'h0f:	  sm4_box_out	<=	8'h05;
		8'h10:	  sm4_box_out	<=	8'h2b;
		8'h11:	  sm4_box_out	<=	8'h67;
		8'h12:	  sm4_box_out	<=	8'h9a;
		8'h13:	  sm4_box_out	<=	8'h76;
		8'h14:	  sm4_box_out	<=	8'h2a;
		8'h15:	  sm4_box_out	<=	8'hbe;
		8'h16:	  sm4_box_out	<=	8'h04;
		8'h17:	  sm4_box_out	<=	8'hc3;
		8'h18:	  sm4_box_out	<=	8'haa;
		8'h19:	  sm4_box_out	<=	8'h44;
		8'h1a:	  sm4_box_out	<=	8'h13;
		8'h1b:	  sm4_box_out	<=	8'h26;
		8'h1c:	  sm4_box_out	<=	8'h49;
		8'h1d:	  sm4_box_out	<=	8'h86;
		8'h1e:	  sm4_box_out	<=	8'h06;
		8'h1f:	  sm4_box_out	<=	8'h99;
		8'h20:	  sm4_box_out	<=	8'h9c;
		8'h21:	  sm4_box_out	<=	8'h42;
		8'h22:	  sm4_box_out	<=	8'h50;
		8'h23:	  sm4_box_out	<=	8'hf4;
		8'h24:	  sm4_box_out	<=	8'h91;
		8'h25:	  sm4_box_out	<=	8'hef;
		8'h26:	  sm4_box_out	<=	8'h98;
		8'h27:	  sm4_box_out	<=	8'h7a;
		8'h28:	  sm4_box_out	<=	8'h33;
		8'h29:	  sm4_box_out	<=	8'h54;
		8'h2a:	  sm4_box_out	<=	8'h0b;
		8'h2b:	  sm4_box_out	<=	8'h43;
		8'h2c:	  sm4_box_out	<=	8'hed;
		8'h2d:	  sm4_box_out	<=	8'hcf;
		8'h2e:	  sm4_box_out	<=	8'hac;
		8'h2f:	  sm4_box_out	<=	8'h62;
		8'h30:	  sm4_box_out	<=	8'he4;
		8'h31:	  sm4_box_out	<=	8'hb3;
		8'h32:	  sm4_box_out	<=	8'h1c;
		8'h33:	  sm4_box_out	<=	8'ha9;
		8'h34:	  sm4_box_out	<=	8'hc9;
		8'h35:	  sm4_box_out	<=	8'h08;
		8'h36:	  sm4_box_out	<=	8'he8;
		8'h37:	  sm4_box_out	<=	8'h95;
		8'h38:	  sm4_box_out	<=	8'h80;
		8'h39:	  sm4_box_out	<=	8'hdf;
		8'h3a:	  sm4_box_out	<=	8'h94;
		8'h3b:	  sm4_box_out	<=	8'hfa;
		8'h3c:	  sm4_box_out	<=	8'h75;
		8'h3d:	  sm4_box_out	<=	8'h8f;
		8'h3e:	  sm4_box_out	<=	8'h3f;
		8'h3f:	  sm4_box_out	<=	8'ha6;
		8'h40:	  sm4_box_out	<=	8'h47;
		8'h41:	  sm4_box_out	<=	8'h07;
		8'h42:	  sm4_box_out	<=	8'ha7;
		8'h43:	  sm4_box_out	<=	8'hfc;
		8'h44:	  sm4_box_out	<=	8'hf3;
		8'h45:	  sm4_box_out	<=	8'h73;
		8'h46:	  sm4_box_out	<=	8'h17;
		8'h47:	  sm4_box_out	<=	8'hba;
		8'h48:	  sm4_box_out	<=	8'h83;
		8'h49:	  sm4_box_out	<=	8'h59;
		8'h4a:	  sm4_box_out	<=	8'h3c;
		8'h4b:	  sm4_box_out	<=	8'h19;
		8'h4c:	  sm4_box_out	<=	8'he6;
		8'h4d:	  sm4_box_out	<=	8'h85;
		8'h4e:	  sm4_box_out	<=	8'h4f;
		8'h4f:	  sm4_box_out	<=	8'ha8;
		8'h50:	  sm4_box_out	<=	8'h68;
		8'h51:	  sm4_box_out	<=	8'h6b;
		8'h52:	  sm4_box_out	<=	8'h81;
		8'h53:	  sm4_box_out	<=	8'hb2;
		8'h54:	  sm4_box_out	<=	8'h71;
		8'h55:	  sm4_box_out	<=	8'h64;
		8'h56:	  sm4_box_out	<=	8'hda;
		8'h57:	  sm4_box_out	<=	8'h8b;
		8'h58:	  sm4_box_out	<=	8'hf8;
		8'h59:	  sm4_box_out	<=	8'heb;
		8'h5a:	  sm4_box_out	<=	8'h0f;
		8'h5b:	  sm4_box_out	<=	8'h4b;
		8'h5c:	  sm4_box_out	<=	8'h70;
		8'h5d:	  sm4_box_out	<=	8'h56;
		8'h5e:	  sm4_box_out	<=	8'h9d;
		8'h5f:	  sm4_box_out	<=	8'h35;
		8'h60:	  sm4_box_out	<=	8'h1e;
		8'h61:	  sm4_box_out	<=	8'h24;
		8'h62:	  sm4_box_out	<=	8'h0e;
		8'h63:	  sm4_box_out	<=	8'h5e;
		8'h64:	  sm4_box_out	<=	8'h63;
		8'h65:	  sm4_box_out	<=	8'h58;
		8'h66:	  sm4_box_out	<=	8'hd1;
		8'h67:	  sm4_box_out	<=	8'ha2;
		8'h68:	  sm4_box_out	<=	8'h25;
		8'h69:	  sm4_box_out	<=	8'h22;
		8'h6a:	  sm4_box_out	<=	8'h7c;
		8'h6b:	  sm4_box_out	<=	8'h3b;
		8'h6c:	  sm4_box_out	<=	8'h01;
		8'h6d:	  sm4_box_out	<=	8'h21;
		8'h6e:	  sm4_box_out	<=	8'h78;
		8'h6f:	  sm4_box_out	<=	8'h87;
		8'h70:	  sm4_box_out	<=	8'hd4;
		8'h71:	  sm4_box_out	<=	8'h00;
		8'h72:	  sm4_box_out	<=	8'h46;
		8'h73:	  sm4_box_out	<=	8'h57;
		8'h74:	  sm4_box_out	<=	8'h9f;
		8'h75:	  sm4_box_out	<=	8'hd3;
		8'h76:	  sm4_box_out	<=	8'h27;
		8'h77:	  sm4_box_out	<=	8'h52;
		8'h78:	  sm4_box_out	<=	8'h4c;
		8'h79:	  sm4_box_out	<=	8'h36;
		8'h7a:	  sm4_box_out	<=	8'h02;
		8'h7b:	  sm4_box_out	<=	8'he7;
		8'h7c:	  sm4_box_out	<=	8'ha0;
		8'h7d:	  sm4_box_out	<=	8'hc4;
		8'h7e:	  sm4_box_out	<=	8'hc8;
		8'h7f:	  sm4_box_out	<=	8'h9e;
		8'h80:	  sm4_box_out	<=	8'hea;
		8'h81:	  sm4_box_out	<=	8'hbf;
		8'h82:	  sm4_box_out	<=	8'h8a;
		8'h83:	  sm4_box_out	<=	8'hd2;
		8'h84:	  sm4_box_out	<=	8'h40;
		8'h85:	  sm4_box_out	<=	8'hc7;
		8'h86:	  sm4_box_out	<=	8'h38;
		8'h87:	  sm4_box_out	<=	8'hb5;
		8'h88:	  sm4_box_out	<=	8'ha3;
		8'h89:	  sm4_box_out	<=	8'hf7;
		8'h8a:	  sm4_box_out	<=	8'hf2;
		8'h8b:	  sm4_box_out	<=	8'hce;
		8'h8c:	  sm4_box_out	<=	8'hf9;
		8'h8d:	  sm4_box_out	<=	8'h61;
		8'h8e:	  sm4_box_out	<=	8'h15;
		8'h8f:	  sm4_box_out	<=	8'ha1;
		8'h90:	  sm4_box_out	<=	8'he0;
		8'h91:	  sm4_box_out	<=	8'hae;
		8'h92:	  sm4_box_out	<=	8'h5d;
		8'h93:	  sm4_box_out	<=	8'ha4;
		8'h94:	  sm4_box_out	<=	8'h9b;
		8'h95:	  sm4_box_out	<=	8'h34;
		8'h96:	  sm4_box_out	<=	8'h1a;
		8'h97:	  sm4_box_out	<=	8'h55;
		8'h98:	  sm4_box_out	<=	8'had;
		8'h99:	  sm4_box_out	<=	8'h93;
		8'h9a:	  sm4_box_out	<=	8'h32;
		8'h9b:	  sm4_box_out	<=	8'h30;
		8'h9c:	  sm4_box_out	<=	8'hf5;
		8'h9d:	  sm4_box_out	<=	8'h8c;
		8'h9e:	  sm4_box_out	<=	8'hb1;
		8'h9f:	  sm4_box_out	<=	8'he3;
		8'ha0:	  sm4_box_out	<=	8'h1d;
		8'ha1:	  sm4_box_out	<=	8'hf6;
		8'ha2:	  sm4_box_out	<=	8'he2;
		8'ha3:	  sm4_box_out	<=	8'h2e;
		8'ha4:	  sm4_box_out	<=	8'h82;
		8'ha5:	  sm4_box_out	<=	8'h66;
		8'ha6:	  sm4_box_out	<=	8'hca;
		8'ha7:	  sm4_box_out	<=	8'h60;
		8'ha8:	  sm4_box_out	<=	8'hc0;
		8'ha9:	  sm4_box_out	<=	8'h29;
		8'haa:	  sm4_box_out	<=	8'h23;
		8'hab:	  sm4_box_out	<=	8'hab;
		8'hac:	  sm4_box_out	<=	8'h0d;
		8'had:	  sm4_box_out	<=	8'h53;
		8'hae:	  sm4_box_out	<=	8'h4e;
		8'haf:	  sm4_box_out	<=	8'h6f;
		8'hb0:	  sm4_box_out	<=	8'hd5;
		8'hb1:	  sm4_box_out	<=	8'hdb;
		8'hb2:	  sm4_box_out	<=	8'h37;
		8'hb3:	  sm4_box_out	<=	8'h45;
		8'hb4:	  sm4_box_out	<=	8'hde;
		8'hb5:	  sm4_box_out	<=	8'hfd;
		8'hb6:	  sm4_box_out	<=	8'h8e;
		8'hb7:	  sm4_box_out	<=	8'h2f;
		8'hb8:	  sm4_box_out	<=	8'h03;
		8'hb9:	  sm4_box_out	<=	8'hff;
		8'hba:	  sm4_box_out	<=	8'h6a;
		8'hbb:	  sm4_box_out	<=	8'h72;
		8'hbc:	  sm4_box_out	<=	8'h6d;
		8'hbd:	  sm4_box_out	<=	8'h6c;
		8'hbe:	  sm4_box_out	<=	8'h5b;
		8'hbf:	  sm4_box_out	<=	8'h51;
		8'hc0:	  sm4_box_out	<=	8'h8d;
		8'hc1:	  sm4_box_out	<=	8'h1b;
		8'hc2:	  sm4_box_out	<=	8'haf;
		8'hc3:	  sm4_box_out	<=	8'h92;
		8'hc4:	  sm4_box_out	<=	8'hbb;
		8'hc5:	  sm4_box_out	<=	8'hdd;
		8'hc6:	  sm4_box_out	<=	8'hbc;
		8'hc7:	  sm4_box_out	<=	8'h7f;
		8'hc8:	  sm4_box_out	<=	8'h11;
		8'hc9:	  sm4_box_out	<=	8'hd9;
		8'hca:	  sm4_box_out	<=	8'h5c;
		8'hcb:	  sm4_box_out	<=	8'h41;
		8'hcc:	  sm4_box_out	<=	8'h1f;
		8'hcd:	  sm4_box_out	<=	8'h10;
		8'hce:	  sm4_box_out	<=	8'h5a;
		8'hcf:	  sm4_box_out	<=	8'hd8;
		8'hd0:	  sm4_box_out	<=	8'h0a;
		8'hd1:	  sm4_box_out	<=	8'hc1;
		8'hd2:	  sm4_box_out	<=	8'h31;
		8'hd3:	  sm4_box_out	<=	8'h88;
		8'hd4:	  sm4_box_out	<=	8'ha5;
		8'hd5:	  sm4_box_out	<=	8'hcd;
		8'hd6:	  sm4_box_out	<=	8'h7b;
		8'hd7:	  sm4_box_out	<=	8'hbd;
		8'hd8:	  sm4_box_out	<=	8'h2d;
		8'hd9:	  sm4_box_out	<=	8'h74;
		8'hda:	  sm4_box_out	<=	8'hd0;
		8'hdb:	  sm4_box_out	<=	8'h12;
		8'hdc:	  sm4_box_out	<=	8'hb8;
		8'hdd:	  sm4_box_out	<=	8'he5;
		8'hde:	  sm4_box_out	<=	8'hb4;
		8'hdf:	  sm4_box_out	<=	8'hb0;
		8'he0:	  sm4_box_out	<=	8'h89;
		8'he1:	  sm4_box_out	<=	8'h69;
		8'he2:	  sm4_box_out	<=	8'h97;
		8'he3:	  sm4_box_out	<=	8'h4a;
		8'he4:	  sm4_box_out	<=	8'h0c;
		8'he5:	  sm4_box_out	<=	8'h96;
		8'he6:	  sm4_box_out	<=	8'h77;
		8'he7:	  sm4_box_out	<=	8'h7e;
		8'he8:	  sm4_box_out	<=	8'h65;
		8'he9:	  sm4_box_out	<=	8'hb9;
		8'hea:	  sm4_box_out	<=	8'hf1;
		8'heb:	  sm4_box_out	<=	8'h09;
		8'hec:	  sm4_box_out	<=	8'hc5;
		8'hed:	  sm4_box_out	<=	8'h6e;
		8'hee:	  sm4_box_out	<=	8'hc6;
		8'hef:	  sm4_box_out	<=	8'h84;
		8'hf0:	  sm4_box_out	<=	8'h18;
		8'hf1:	  sm4_box_out	<=	8'hf0;
		8'hf2:	  sm4_box_out	<=	8'h7d;
		8'hf3:	  sm4_box_out	<=	8'hec;
		8'hf4:	  sm4_box_out	<=	8'h3a;
		8'hf5:	  sm4_box_out	<=	8'hdc;
		8'hf6:	  sm4_box_out	<=	8'h4d;
		8'hf7:	  sm4_box_out	<=	8'h20;
		8'hf8:	  sm4_box_out	<=	8'h79;
		8'hf9:	  sm4_box_out	<=	8'hee;
		8'hfa:	  sm4_box_out	<=	8'h5f;
		8'hfb:	  sm4_box_out	<=	8'h3e;
		8'hfc:	  sm4_box_out	<=	8'hd7;
		8'hfd:	  sm4_box_out	<=	8'hcb;
		8'hfe:	  sm4_box_out	<=	8'h39;
		default:  sm4_box_out	<=	8'h48; //8'hff
	endcase
end

endmodule
